`include "ethernet_frame_pkg.sv"
`include "axi_master_model.sv"
`include "axi_slave_model.sv"
`include "eth_tx_protocol_check.sv"
`include "AXI_interface.sv"
`include "rtl_struct.sv"
`include "eth_core.sv"
`include "eth_tx.sv"
`include "dma_controller_tx.sv"
`include "AXI_master.sv"
`include "AXI_slave.sv"
`include "CRC32_D8.sv"
`include "CRC32_D16.sv"
`include "CRC32_D24.sv"
`include "CRC32_D32.sv"
`include "CRC32_D40.sv"
`include "CRC32_D48.sv"
`include "CRC32_D56.sv"
`include "CRC32_D64.sv"
`include "CRC_block.sv"
`include "eth_tx_crc.sv"
`include "dma_fifo.sv"
`include "rs_layer.sv"
`include "prienc.sv"
`include "QOS_arb.sv"
`include "queue_selection.sv"
//`include "dma_fifo_exmem.sv"
`include "dma_fifo_exmem_crc.sv"
`include "dma_fifo_exmem_pktd.sv"
`include "dma_fifo_exmem_pktc.sv"
`include "dma_fifo_exmem_swchaddr.sv"
`include "dma_fifo_exmem_swchdata.sv"
`include "dma_fifo_exmem_swchrsp.sv"
//`include "mem_model.sv"
`include "mem_model_crc.sv"
`include "mem_model_pktd.sv"
`include "mem_model_pktc.sv"
`include "mem_model_swchaddr.sv"
`include "mem_model_swchdata.sv"
`include "mem_model_swchrsp.sv"
